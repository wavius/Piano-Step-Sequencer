// Adapted fromm Audio_Controller.v

module DAC_controller (
		// Host side
		CLOCK_50,
		reset,
		audio_in_signed,
		//	I2C Side
		DAC_I2C_SCLK,
		DAC_I2C_SDAT	
);
	// Host Side
	input		 		CLOCK_50;
	input		 		reset;
	input signed [31:0] audio_in_signed;
	// I2C Side
	output		 		DAC_I2C_SCLK;
	inout		 		DAC_I2C_SDAT;
	// Internal Registers/Wires
	reg	[15:0]	 		mI2C_CLK_DIV;
	reg	[31:0]	 		mI2C_DATA;
	reg			 		mI2C_CTRL_CLK;
	reg			 		mI2C_GO;
	wire		 		mI2C_END;
	wire		 		mI2C_ACK;
	wire		 		iRST_N 			  = !reset;

	wire [31:0] 		audio_in_unsigned = audio_in_signed + 31'h7FFFFFFF; // shift audio_in to unsigned range
	wire [11:0] 		audio_in_12b      = audio_in_unsigned[31:20];       // audio_in_unsigned / 16

	// Clock Setting
	parameter CLK_Freq		= 50_000_000;  // 50  MHz
	parameter I2C_Freq		= 400_000;	   // 400 KHz

	// I2C
	parameter SLAVE_ADDR    = 8'b11000000; // MCP4625A1T
	parameter CMD_WRITE_DAC = 8'b01000000;

	// Sequential Logic
	// I2C control clock
	always@(posedge CLOCK_50 or negedge iRST_N)
	begin
		if(!iRST_N)
		begin
			mI2C_CTRL_CLK <= 0;
			mI2C_CLK_DIV  <= 0;
		end
		else
		begin
			if( mI2C_CLK_DIV	< (CLK_Freq/I2C_Freq) )
				mI2C_CLK_DIV  <= mI2C_CLK_DIV+1;
			else
			begin
				mI2C_CLK_DIV  <= 0;
				mI2C_CTRL_CLK <= ~mI2C_CTRL_CLK;
			end
		end
	end

	// I2C data driver
	always@(posedge mI2C_CTRL_CLK or negedge iRST_N)
	begin
		if (!iRST_N)
		begin
			mI2C_DATA <= 0;
			mI2C_GO	  <= 0;
		end
		else
		if (!mI2C_GO && mI2C_END)
		begin
			mI2C_DATA <= {SLAVE_ADDR, CMD_WRITE_DAC, audio_in_12b[11:4], {audio_in_12b[3:0], 4'b0000}};
			mI2C_GO   <= 1;
		end
		else if (mI2C_END)
		begin
			mI2C_GO   <= 0;
		end
	end

	// Internal modules
	I2C_Controller_DAC 	U1	(	
			.CLOCK(mI2C_CTRL_CLK),			//	Controller Work Clock
			.DAC_I2C_SCLK(DAC_I2C_SCLK),    //	I2C CLOCK
			.DAC_I2C_SDAT(DAC_I2C_SDAT),	//	I2C DATA
			.I2C_DATA(mI2C_DATA),			//  DATA:[SLAVE_ADDR, CMD, DATA_MSB, DATA_LSB]
			.GO(mI2C_GO),      				//	GO transfor
			.END(mI2C_END),					//	END transfor 
			.ACK(mI2C_ACK),					//	ACK
			.RESET(iRST_N)	
	);

endmodule
