module rom256x16 (
    input [7:0] address,
    input clock,
    output reg [15:0] q
);
    reg [15:0] mem [0:255];
    initial $readmemh("sine256.hex", mem);

    always @(posedge clock)
        q <= mem[address];
endmodule